// instruction fetch unit
`include "define/const.v"
`include "define/inst.v"

module ifu (
    input wire clk, input wire rst
  );
endmodule
