`ifndef UTIL_DFF_V
`define UTIL_DFF_V

module dff #(
    parameter width = 32
  )(
    input wire clk, input wire rst,
    input wire[width - 1: 0] d, output reg[width - 1: 0] q
  );

  always @ (posedge clk or posedge rst) begin
    if (rst) begin
      q <= 0;
    end
    else begin
      q <= d;
    end
  end

endmodule

`endif